module main

// TODO: To be implemented!
